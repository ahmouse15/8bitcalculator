module test (
	input [3:0] in,
	output reg [6:0] out
	);
	
endmodule
