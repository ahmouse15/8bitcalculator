module signed_bcd2bin();

endmodule
