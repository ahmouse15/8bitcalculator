module main();
	input_unit();
endmodule
